
module NIOS_II_Core (
	clk_clk,
	leds_export);	

	input		clk_clk;
	output	[1:0]	leds_export;
endmodule
